package const_float;
parameter float_exp_width = 8;
parameter float_mant_width = 23;
parameter float_width = float_exp_width + float_mant_width + 1;
endpackage 
