package mem_small;
parameter mem_simulated_delay = 5;
parameter memory_size = 16;
endpackage